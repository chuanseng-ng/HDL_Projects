`define ADDR_WIDTH 32
`define DATA_WIDTH 16
`define INSTR_NUM  15
`define ALU_SIZE   8
`define SHIFT_BIT  1
`define MEM_SIZE   256
