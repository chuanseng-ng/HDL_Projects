`ifndef FIFO_MEM_REGS_PKG__SV
`define FIFO_MEM_REGS_PKG__SV

  package fifo_mem_regs_pkg;

    // Import UVM
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Include Reg Model UVCs

  endpackage

`endif

//End of fifo_mem_regs_pkg
